// Copyright (c) 2020 Stunx (Jose Mendoza). All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module scanner


