// Copyright (c) 2020 StunxFS. All rights reserved. Use of this source code is
// governed by an MIT license that can be found in the LICENSE file.
module about

pub const (
	version 			= "0.1.0a0"
	gen_bin_version 	= "alpha0" // Más tarde: 0.1.0a
	build_time			= '<unknown>'
)

