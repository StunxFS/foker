// Copyright (c) 2020 Stunx. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module about

pub const (
	version = "0.1.0.alpha.0"
)

